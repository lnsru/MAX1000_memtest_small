-- NIOS_test_board.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity NIOS_test_board is
	port (
		clk_in_clk      : in    std_logic                     := '0';             --    clk_in.clk
		pio_led_export  : out   std_logic_vector(7 downto 0);                     --   pio_led.export
		pio_mode_export : in    std_logic_vector(2 downto 0)  := (others => '0'); --  pio_mode.export
		reset_reset_n   : in    std_logic                     := '0';             --     reset.reset_n
		sdram_addr      : out   std_logic_vector(11 downto 0);                    --     sdram.addr
		sdram_ba        : out   std_logic_vector(1 downto 0);                     --          .ba
		sdram_cas_n     : out   std_logic;                                        --          .cas_n
		sdram_cke       : out   std_logic;                                        --          .cke
		sdram_cs_n      : out   std_logic;                                        --          .cs_n
		sdram_dq        : inout std_logic_vector(15 downto 0) := (others => '0'); --          .dq
		sdram_dqm       : out   std_logic_vector(1 downto 0);                     --          .dqm
		sdram_ras_n     : out   std_logic;                                        --          .ras_n
		sdram_we_n      : out   std_logic;                                        --          .we_n
		sdram_clk_clk   : out   std_logic;                                        -- sdram_clk.clk
		spi_flash_MISO  : in    std_logic                     := '0';             -- spi_flash.MISO
		spi_flash_MOSI  : out   std_logic;                                        --          .MOSI
		spi_flash_SCLK  : out   std_logic;                                        --          .SCLK
		spi_flash_SS_n  : out   std_logic;                                        --          .SS_n
		spi_g_sen_MISO  : in    std_logic                     := '0';             -- spi_g_sen.MISO
		spi_g_sen_MOSI  : out   std_logic;                                        --          .MOSI
		spi_g_sen_SCLK  : out   std_logic;                                        --          .SCLK
		spi_g_sen_SS_n  : out   std_logic;                                        --          .SS_n
		uart_rxd        : in    std_logic                     := '0';             --      uart.rxd
		uart_txd        : out   std_logic                                         --          .txd
	);
end entity NIOS_test_board;

architecture rtl of NIOS_test_board is
	component NIOS_test_board_nios2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(24 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component NIOS_test_board_nios2;

	component altera_onchip_flash is
		generic (
			INIT_FILENAME                       : string  := "";
			INIT_FILENAME_SIM                   : string  := "";
			DEVICE_FAMILY                       : string  := "Unknown";
			PART_NAME                           : string  := "Unknown";
			DEVICE_ID                           : string  := "Unknown";
			SECTOR1_START_ADDR                  : integer := 0;
			SECTOR1_END_ADDR                    : integer := 0;
			SECTOR2_START_ADDR                  : integer := 0;
			SECTOR2_END_ADDR                    : integer := 0;
			SECTOR3_START_ADDR                  : integer := 0;
			SECTOR3_END_ADDR                    : integer := 0;
			SECTOR4_START_ADDR                  : integer := 0;
			SECTOR4_END_ADDR                    : integer := 0;
			SECTOR5_START_ADDR                  : integer := 0;
			SECTOR5_END_ADDR                    : integer := 0;
			MIN_VALID_ADDR                      : integer := 0;
			MAX_VALID_ADDR                      : integer := 0;
			MIN_UFM_VALID_ADDR                  : integer := 0;
			MAX_UFM_VALID_ADDR                  : integer := 0;
			SECTOR1_MAP                         : integer := 0;
			SECTOR2_MAP                         : integer := 0;
			SECTOR3_MAP                         : integer := 0;
			SECTOR4_MAP                         : integer := 0;
			SECTOR5_MAP                         : integer := 0;
			ADDR_RANGE1_END_ADDR                : integer := 0;
			ADDR_RANGE2_END_ADDR                : integer := 0;
			ADDR_RANGE1_OFFSET                  : integer := 0;
			ADDR_RANGE2_OFFSET                  : integer := 0;
			ADDR_RANGE3_OFFSET                  : integer := 0;
			AVMM_DATA_ADDR_WIDTH                : integer := 19;
			AVMM_DATA_DATA_WIDTH                : integer := 32;
			AVMM_DATA_BURSTCOUNT_WIDTH          : integer := 4;
			SECTOR_READ_PROTECTION_MODE         : integer := 31;
			FLASH_SEQ_READ_DATA_COUNT           : integer := 2;
			FLASH_ADDR_ALIGNMENT_BITS           : integer := 1;
			FLASH_READ_CYCLE_MAX_INDEX          : integer := 4;
			FLASH_RESET_CYCLE_MAX_INDEX         : integer := 29;
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  : integer := 112;
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX : integer := 40603248;
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX : integer := 35382;
			PARALLEL_MODE                       : boolean := true;
			READ_AND_WRITE_MODE                 : boolean := true;
			WRAPPING_BURST_MODE                 : boolean := false;
			IS_DUAL_BOOT                        : string  := "False";
			IS_ERAM_SKIP                        : string  := "False";
			IS_COMPRESSED_IMAGE                 : string  := "False"
		);
		port (
			clock                   : in  std_logic                     := 'X';             -- clk
			reset_n                 : in  std_logic                     := 'X';             -- reset_n
			avmm_data_addr          : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			avmm_data_read          : in  std_logic                     := 'X';             -- read
			avmm_data_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_data_write         : in  std_logic                     := 'X';             -- write
			avmm_data_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_data_waitrequest   : out std_logic;                                        -- waitrequest
			avmm_data_readdatavalid : out std_logic;                                        -- readdatavalid
			avmm_data_burstcount    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			avmm_csr_addr           : in  std_logic                     := 'X';             -- address
			avmm_csr_read           : in  std_logic                     := 'X';             -- read
			avmm_csr_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_csr_write          : in  std_logic                     := 'X';             -- write
			avmm_csr_readdata       : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component altera_onchip_flash;

	component NIOS_test_board_onchip_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component NIOS_test_board_onchip_ram;

	component NIOS_test_board_pio_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component NIOS_test_board_pio_led;

	component NIOS_test_board_pio_mode is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- export
		);
	end component NIOS_test_board_pio_mode;

	component NIOS_test_board_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component NIOS_test_board_pll;

	component NIOS_test_board_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component NIOS_test_board_sdram_controller;

	component NIOS_test_board_spi_flash is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component NIOS_test_board_spi_flash;

	component NIOS_test_board_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component NIOS_test_board_sysid;

	component NIOS_test_board_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component NIOS_test_board_uart;

	component NIOS_test_board_mm_interconnect_0 is
		port (
			clk_clk_clk                                           : in  std_logic                     := 'X';             -- clk
			pll_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			nios2_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_data_master_address                             : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			nios2_data_master_waitrequest                         : out std_logic;                                        -- waitrequest
			nios2_data_master_byteenable                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_data_master_read                                : in  std_logic                     := 'X';             -- read
			nios2_data_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_data_master_write                               : in  std_logic                     := 'X';             -- write
			nios2_data_master_writedata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_data_master_debugaccess                         : in  std_logic                     := 'X';             -- debugaccess
			nios2_instruction_master_address                      : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			nios2_instruction_master_waitrequest                  : out std_logic;                                        -- waitrequest
			nios2_instruction_master_read                         : in  std_logic                     := 'X';             -- read
			nios2_instruction_master_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_debug_mem_slave_address                         : out std_logic_vector(8 downto 0);                     -- address
			nios2_debug_mem_slave_write                           : out std_logic;                                        -- write
			nios2_debug_mem_slave_read                            : out std_logic;                                        -- read
			nios2_debug_mem_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_debug_mem_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_debug_mem_slave_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_debug_mem_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			nios2_debug_mem_slave_debugaccess                     : out std_logic;                                        -- debugaccess
			onchip_flash_csr_address                              : out std_logic_vector(0 downto 0);                     -- address
			onchip_flash_csr_write                                : out std_logic;                                        -- write
			onchip_flash_csr_read                                 : out std_logic;                                        -- read
			onchip_flash_csr_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_csr_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_data_address                             : out std_logic_vector(16 downto 0);                    -- address
			onchip_flash_data_write                               : out std_logic;                                        -- write
			onchip_flash_data_read                                : out std_logic;                                        -- read
			onchip_flash_data_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_data_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_data_burstcount                          : out std_logic_vector(3 downto 0);                     -- burstcount
			onchip_flash_data_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			onchip_flash_data_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			onchip_ram_s1_address                                 : out std_logic_vector(12 downto 0);                    -- address
			onchip_ram_s1_write                                   : out std_logic;                                        -- write
			onchip_ram_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                                   : out std_logic;                                        -- clken
			pio_led_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			pio_led_s1_write                                      : out std_logic;                                        -- write
			pio_led_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_led_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			pio_led_s1_chipselect                                 : out std_logic;                                        -- chipselect
			pio_mode_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			pio_mode_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pll_pll_slave_write                                   : out std_logic;                                        -- write
			pll_pll_slave_read                                    : out std_logic;                                        -- read
			pll_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_controller_s1_address                           : out std_logic_vector(21 downto 0);                    -- address
			sdram_controller_s1_write                             : out std_logic;                                        -- write
			sdram_controller_s1_read                              : out std_logic;                                        -- read
			sdram_controller_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                        : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                        : out std_logic;                                        -- chipselect
			spi_flash_spi_control_port_address                    : out std_logic_vector(2 downto 0);                     -- address
			spi_flash_spi_control_port_write                      : out std_logic;                                        -- write
			spi_flash_spi_control_port_read                       : out std_logic;                                        -- read
			spi_flash_spi_control_port_readdata                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_flash_spi_control_port_writedata                  : out std_logic_vector(15 downto 0);                    -- writedata
			spi_flash_spi_control_port_chipselect                 : out std_logic;                                        -- chipselect
			spi_g_sensor_spi_control_port_address                 : out std_logic_vector(2 downto 0);                     -- address
			spi_g_sensor_spi_control_port_write                   : out std_logic;                                        -- write
			spi_g_sensor_spi_control_port_read                    : out std_logic;                                        -- read
			spi_g_sensor_spi_control_port_readdata                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_g_sensor_spi_control_port_writedata               : out std_logic_vector(15 downto 0);                    -- writedata
			spi_g_sensor_spi_control_port_chipselect              : out std_logic;                                        -- chipselect
			sysid_control_slave_address                           : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uart_s1_address                                       : out std_logic_vector(2 downto 0);                     -- address
			uart_s1_write                                         : out std_logic;                                        -- write
			uart_s1_read                                          : out std_logic;                                        -- read
			uart_s1_readdata                                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_s1_writedata                                     : out std_logic_vector(15 downto 0);                    -- writedata
			uart_s1_begintransfer                                 : out std_logic;                                        -- begintransfer
			uart_s1_chipselect                                    : out std_logic                                         -- chipselect
		);
	end component NIOS_test_board_mm_interconnect_0;

	component NIOS_test_board_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component NIOS_test_board_irq_mapper;

	component nios_test_board_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_test_board_rst_controller;

	component nios_test_board_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios_test_board_rst_controller_001;

	signal pll_c0_clk                                                      : std_logic;                     -- pll:c0 -> [irq_mapper:clk, mm_interconnect_0:pll_c0_clk, nios2:clk, onchip_flash:clock, onchip_ram:clk, pio_led:clk, pio_mode:clk, rst_controller:clk, sdram_controller:clk, spi_flash:clk, spi_g_sensor:clk, sysid:clock, uart:clk]
	signal nios2_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	signal nios2_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	signal nios2_data_master_debugaccess                                   : std_logic;                     -- nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	signal nios2_data_master_address                                       : std_logic_vector(24 downto 0); -- nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	signal nios2_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	signal nios2_data_master_read                                          : std_logic;                     -- nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	signal nios2_data_master_write                                         : std_logic;                     -- nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	signal nios2_data_master_writedata                                     : std_logic_vector(31 downto 0); -- nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	signal nios2_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	signal nios2_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	signal nios2_instruction_master_address                                : std_logic_vector(24 downto 0); -- nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	signal nios2_instruction_master_read                                   : std_logic;                     -- nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	signal mm_interconnect_0_sysid_control_slave_readdata                  : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                   : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_onchip_flash_csr_readdata                     : std_logic_vector(31 downto 0); -- onchip_flash:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_csr_readdata
	signal mm_interconnect_0_onchip_flash_csr_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:onchip_flash_csr_address -> onchip_flash:avmm_csr_addr
	signal mm_interconnect_0_onchip_flash_csr_read                         : std_logic;                     -- mm_interconnect_0:onchip_flash_csr_read -> onchip_flash:avmm_csr_read
	signal mm_interconnect_0_onchip_flash_csr_write                        : std_logic;                     -- mm_interconnect_0:onchip_flash_csr_write -> onchip_flash:avmm_csr_write
	signal mm_interconnect_0_onchip_flash_csr_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_flash_csr_writedata -> onchip_flash:avmm_csr_writedata
	signal mm_interconnect_0_onchip_flash_data_readdata                    : std_logic_vector(31 downto 0); -- onchip_flash:avmm_data_readdata -> mm_interconnect_0:onchip_flash_data_readdata
	signal mm_interconnect_0_onchip_flash_data_waitrequest                 : std_logic;                     -- onchip_flash:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_data_waitrequest
	signal mm_interconnect_0_onchip_flash_data_address                     : std_logic_vector(16 downto 0); -- mm_interconnect_0:onchip_flash_data_address -> onchip_flash:avmm_data_addr
	signal mm_interconnect_0_onchip_flash_data_read                        : std_logic;                     -- mm_interconnect_0:onchip_flash_data_read -> onchip_flash:avmm_data_read
	signal mm_interconnect_0_onchip_flash_data_readdatavalid               : std_logic;                     -- onchip_flash:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_data_readdatavalid
	signal mm_interconnect_0_onchip_flash_data_write                       : std_logic;                     -- mm_interconnect_0:onchip_flash_data_write -> onchip_flash:avmm_data_write
	signal mm_interconnect_0_onchip_flash_data_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_flash_data_writedata -> onchip_flash:avmm_data_writedata
	signal mm_interconnect_0_onchip_flash_data_burstcount                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_flash_data_burstcount -> onchip_flash:avmm_data_burstcount
	signal mm_interconnect_0_nios2_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_debug_mem_slave_waitrequest             : std_logic;                     -- nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	signal mm_interconnect_0_nios2_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	signal mm_interconnect_0_nios2_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	signal mm_interconnect_0_nios2_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	signal mm_interconnect_0_pll_pll_slave_readdata                        : std_logic_vector(31 downto 0); -- pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	signal mm_interconnect_0_pll_pll_slave_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pll_pll_slave_address -> pll:address
	signal mm_interconnect_0_pll_pll_slave_read                            : std_logic;                     -- mm_interconnect_0:pll_pll_slave_read -> pll:read
	signal mm_interconnect_0_pll_pll_slave_write                           : std_logic;                     -- mm_interconnect_0:pll_pll_slave_write -> pll:write
	signal mm_interconnect_0_pll_pll_slave_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	signal mm_interconnect_0_onchip_ram_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata                        : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address                         : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal mm_interconnect_0_sdram_controller_s1_chipselect                : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                  : std_logic_vector(15 downto 0); -- sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest               : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                   : std_logic_vector(21 downto 0); -- mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                      : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid             : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                     : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal mm_interconnect_0_pio_led_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	signal mm_interconnect_0_pio_led_s1_readdata                           : std_logic_vector(31 downto 0); -- pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	signal mm_interconnect_0_pio_led_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_led_s1_address -> pio_led:address
	signal mm_interconnect_0_pio_led_s1_write                              : std_logic;                     -- mm_interconnect_0:pio_led_s1_write -> mm_interconnect_0_pio_led_s1_write:in
	signal mm_interconnect_0_pio_led_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	signal mm_interconnect_0_uart_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	signal mm_interconnect_0_uart_s1_readdata                              : std_logic_vector(15 downto 0); -- uart:readdata -> mm_interconnect_0:uart_s1_readdata
	signal mm_interconnect_0_uart_s1_address                               : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_s1_address -> uart:address
	signal mm_interconnect_0_uart_s1_read                                  : std_logic;                     -- mm_interconnect_0:uart_s1_read -> mm_interconnect_0_uart_s1_read:in
	signal mm_interconnect_0_uart_s1_begintransfer                         : std_logic;                     -- mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	signal mm_interconnect_0_uart_s1_write                                 : std_logic;                     -- mm_interconnect_0:uart_s1_write -> mm_interconnect_0_uart_s1_write:in
	signal mm_interconnect_0_uart_s1_writedata                             : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_s1_writedata -> uart:writedata
	signal mm_interconnect_0_pio_mode_s1_readdata                          : std_logic_vector(31 downto 0); -- pio_mode:readdata -> mm_interconnect_0:pio_mode_s1_readdata
	signal mm_interconnect_0_pio_mode_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_mode_s1_address -> pio_mode:address
	signal mm_interconnect_0_spi_flash_spi_control_port_chipselect         : std_logic;                     -- mm_interconnect_0:spi_flash_spi_control_port_chipselect -> spi_flash:spi_select
	signal mm_interconnect_0_spi_flash_spi_control_port_readdata           : std_logic_vector(15 downto 0); -- spi_flash:data_to_cpu -> mm_interconnect_0:spi_flash_spi_control_port_readdata
	signal mm_interconnect_0_spi_flash_spi_control_port_address            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_flash_spi_control_port_address -> spi_flash:mem_addr
	signal mm_interconnect_0_spi_flash_spi_control_port_read               : std_logic;                     -- mm_interconnect_0:spi_flash_spi_control_port_read -> mm_interconnect_0_spi_flash_spi_control_port_read:in
	signal mm_interconnect_0_spi_flash_spi_control_port_write              : std_logic;                     -- mm_interconnect_0:spi_flash_spi_control_port_write -> mm_interconnect_0_spi_flash_spi_control_port_write:in
	signal mm_interconnect_0_spi_flash_spi_control_port_writedata          : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_flash_spi_control_port_writedata -> spi_flash:data_from_cpu
	signal mm_interconnect_0_spi_g_sensor_spi_control_port_chipselect      : std_logic;                     -- mm_interconnect_0:spi_g_sensor_spi_control_port_chipselect -> spi_g_sensor:spi_select
	signal mm_interconnect_0_spi_g_sensor_spi_control_port_readdata        : std_logic_vector(15 downto 0); -- spi_g_sensor:data_to_cpu -> mm_interconnect_0:spi_g_sensor_spi_control_port_readdata
	signal mm_interconnect_0_spi_g_sensor_spi_control_port_address         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_g_sensor_spi_control_port_address -> spi_g_sensor:mem_addr
	signal mm_interconnect_0_spi_g_sensor_spi_control_port_read            : std_logic;                     -- mm_interconnect_0:spi_g_sensor_spi_control_port_read -> mm_interconnect_0_spi_g_sensor_spi_control_port_read:in
	signal mm_interconnect_0_spi_g_sensor_spi_control_port_write           : std_logic;                     -- mm_interconnect_0:spi_g_sensor_spi_control_port_write -> mm_interconnect_0_spi_g_sensor_spi_control_port_write:in
	signal mm_interconnect_0_spi_g_sensor_spi_control_port_writedata       : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_g_sensor_spi_control_port_writedata -> spi_g_sensor:data_from_cpu
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- uart:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- spi_flash:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- spi_g_sensor:irq -> irq_mapper:receiver2_irq
	signal nios2_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, onchip_ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [nios2:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	signal nios2_debug_reset_request_reset                                 : std_logic;                     -- nios2:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv            : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv      : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal mm_interconnect_0_pio_led_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_pio_led_s1_write:inv -> pio_led:write_n
	signal mm_interconnect_0_uart_s1_read_ports_inv                        : std_logic;                     -- mm_interconnect_0_uart_s1_read:inv -> uart:read_n
	signal mm_interconnect_0_uart_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_uart_s1_write:inv -> uart:write_n
	signal mm_interconnect_0_spi_flash_spi_control_port_read_ports_inv     : std_logic;                     -- mm_interconnect_0_spi_flash_spi_control_port_read:inv -> spi_flash:read_n
	signal mm_interconnect_0_spi_flash_spi_control_port_write_ports_inv    : std_logic;                     -- mm_interconnect_0_spi_flash_spi_control_port_write:inv -> spi_flash:write_n
	signal mm_interconnect_0_spi_g_sensor_spi_control_port_read_ports_inv  : std_logic;                     -- mm_interconnect_0_spi_g_sensor_spi_control_port_read:inv -> spi_g_sensor:read_n
	signal mm_interconnect_0_spi_g_sensor_spi_control_port_write_ports_inv : std_logic;                     -- mm_interconnect_0_spi_g_sensor_spi_control_port_write:inv -> spi_g_sensor:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [nios2:reset_n, onchip_flash:reset_n, pio_led:reset_n, pio_mode:reset_n, sdram_controller:reset_n, spi_flash:reset_n, spi_g_sensor:reset_n, sysid:reset_n, uart:reset_n]

begin

	nios2 : component NIOS_test_board_nios2
		port map (
			clk                                 => pll_c0_clk,                                          --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => nios2_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_data_master_read,                              --                          .read
			d_readdata                          => nios2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_data_master_write,                             --                          .write
			d_writedata                         => nios2_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	onchip_flash : component altera_onchip_flash
		generic map (
			INIT_FILENAME                       => "",
			INIT_FILENAME_SIM                   => "",
			DEVICE_FAMILY                       => "MAX 10",
			PART_NAME                           => "10M08SAU169C8G",
			DEVICE_ID                           => "08",
			SECTOR1_START_ADDR                  => 0,
			SECTOR1_END_ADDR                    => 4095,
			SECTOR2_START_ADDR                  => 4096,
			SECTOR2_END_ADDR                    => 8191,
			SECTOR3_START_ADDR                  => 8192,
			SECTOR3_END_ADDR                    => 29183,
			SECTOR4_START_ADDR                  => 29184,
			SECTOR4_END_ADDR                    => 44031,
			SECTOR5_START_ADDR                  => 44032,
			SECTOR5_END_ADDR                    => 79871,
			MIN_VALID_ADDR                      => 0,
			MAX_VALID_ADDR                      => 79871,
			MIN_UFM_VALID_ADDR                  => 0,
			MAX_UFM_VALID_ADDR                  => 8191,
			SECTOR1_MAP                         => 1,
			SECTOR2_MAP                         => 2,
			SECTOR3_MAP                         => 3,
			SECTOR4_MAP                         => 4,
			SECTOR5_MAP                         => 5,
			ADDR_RANGE1_END_ADDR                => 79871,
			ADDR_RANGE2_END_ADDR                => 79871,
			ADDR_RANGE1_OFFSET                  => 512,
			ADDR_RANGE2_OFFSET                  => 0,
			ADDR_RANGE3_OFFSET                  => 0,
			AVMM_DATA_ADDR_WIDTH                => 17,
			AVMM_DATA_DATA_WIDTH                => 32,
			AVMM_DATA_BURSTCOUNT_WIDTH          => 4,
			SECTOR_READ_PROTECTION_MODE         => 0,
			FLASH_SEQ_READ_DATA_COUNT           => 2,
			FLASH_ADDR_ALIGNMENT_BITS           => 1,
			FLASH_READ_CYCLE_MAX_INDEX          => 4,
			FLASH_RESET_CYCLE_MAX_INDEX         => 12,
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  => 60,
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX => 17500000,
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX => 15250,
			PARALLEL_MODE                       => true,
			READ_AND_WRITE_MODE                 => true,
			WRAPPING_BURST_MODE                 => false,
			IS_DUAL_BOOT                        => "False",
			IS_ERAM_SKIP                        => "False",
			IS_COMPRESSED_IMAGE                 => "False"
		)
		port map (
			clock                   => pll_c0_clk,                                        --    clk.clk
			reset_n                 => rst_controller_reset_out_reset_ports_inv,          -- nreset.reset_n
			avmm_data_addr          => mm_interconnect_0_onchip_flash_data_address,       --   data.address
			avmm_data_read          => mm_interconnect_0_onchip_flash_data_read,          --       .read
			avmm_data_writedata     => mm_interconnect_0_onchip_flash_data_writedata,     --       .writedata
			avmm_data_write         => mm_interconnect_0_onchip_flash_data_write,         --       .write
			avmm_data_readdata      => mm_interconnect_0_onchip_flash_data_readdata,      --       .readdata
			avmm_data_waitrequest   => mm_interconnect_0_onchip_flash_data_waitrequest,   --       .waitrequest
			avmm_data_readdatavalid => mm_interconnect_0_onchip_flash_data_readdatavalid, --       .readdatavalid
			avmm_data_burstcount    => mm_interconnect_0_onchip_flash_data_burstcount,    --       .burstcount
			avmm_csr_addr           => mm_interconnect_0_onchip_flash_csr_address(0),     --    csr.address
			avmm_csr_read           => mm_interconnect_0_onchip_flash_csr_read,           --       .read
			avmm_csr_writedata      => mm_interconnect_0_onchip_flash_csr_writedata,      --       .writedata
			avmm_csr_write          => mm_interconnect_0_onchip_flash_csr_write,          --       .write
			avmm_csr_readdata       => mm_interconnect_0_onchip_flash_csr_readdata        --       .readdata
		);

	onchip_ram : component NIOS_test_board_onchip_ram
		port map (
			clk        => pll_c0_clk,                                 --   clk1.clk
			address    => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	pio_led : component NIOS_test_board_pio_led
		port map (
			clk        => pll_c0_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_pio_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_led_s1_readdata,        --                    .readdata
			out_port   => pio_led_export                                -- external_connection.export
		);

	pio_mode : component NIOS_test_board_pio_mode
		port map (
			clk      => pll_c0_clk,                               --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_pio_mode_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_pio_mode_s1_readdata,   --                    .readdata
			in_port  => pio_mode_export                           -- external_connection.export
		);

	pll : component NIOS_test_board_pll
		port map (
			clk                => clk_in_clk,                                --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,        -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_pll_slave_writedata, --                      .writedata
			c0                 => pll_c0_clk,                                --                    c0.clk
			c1                 => sdram_clk_clk,                             --                    c1.clk
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			c2                 => open,                                      --           (terminated)
			c3                 => open,                                      --           (terminated)
			c4                 => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			locked             => open,                                      --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "000",                                     --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	sdram_controller : component NIOS_test_board_sdram_controller
		port map (
			clk            => pll_c0_clk,                                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                   -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                                 --  wire.export
			zs_ba          => sdram_ba,                                                   --      .export
			zs_cas_n       => sdram_cas_n,                                                --      .export
			zs_cke         => sdram_cke,                                                  --      .export
			zs_cs_n        => sdram_cs_n,                                                 --      .export
			zs_dq          => sdram_dq,                                                   --      .export
			zs_dqm         => sdram_dqm,                                                  --      .export
			zs_ras_n       => sdram_ras_n,                                                --      .export
			zs_we_n        => sdram_we_n                                                  --      .export
		);

	spi_flash : component NIOS_test_board_spi_flash
		port map (
			clk           => pll_c0_clk,                                                   --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                     --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_flash_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_flash_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_flash_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_flash_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_flash_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_flash_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver1_irq,                                     --              irq.irq
			MISO          => spi_flash_MISO,                                               --         external.export
			MOSI          => spi_flash_MOSI,                                               --                 .export
			SCLK          => spi_flash_SCLK,                                               --                 .export
			SS_n          => spi_flash_SS_n                                                --                 .export
		);

	spi_g_sensor : component NIOS_test_board_spi_flash
		port map (
			clk           => pll_c0_clk,                                                      --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                        --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_g_sensor_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_g_sensor_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_g_sensor_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_g_sensor_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_g_sensor_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_g_sensor_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver2_irq,                                        --              irq.irq
			MISO          => spi_g_sen_MISO,                                                  --         external.export
			MOSI          => spi_g_sen_MOSI,                                                  --                 .export
			SCLK          => spi_g_sen_SCLK,                                                  --                 .export
			SS_n          => spi_g_sen_SS_n                                                   --                 .export
		);

	sysid : component NIOS_test_board_sysid
		port map (
			clock    => pll_c0_clk,                                       --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	uart : component NIOS_test_board_uart
		port map (
			clk           => pll_c0_clk,                                --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address       => mm_interconnect_0_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_s1_readdata,        --                    .readdata
			rxd           => uart_rxd,                                  -- external_connection.export
			txd           => uart_txd,                                  --                    .export
			irq           => irq_mapper_receiver0_irq                   --                 irq.irq
		);

	mm_interconnect_0 : component NIOS_test_board_mm_interconnect_0
		port map (
			clk_clk_clk                                           => clk_in_clk,                                                 --                                         clk_clk.clk
			pll_c0_clk                                            => pll_c0_clk,                                                 --                                          pll_c0.clk
			nios2_reset_reset_bridge_in_reset_reset               => rst_controller_reset_out_reset,                             --               nios2_reset_reset_bridge_in_reset.reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                         -- pll_inclk_interface_reset_reset_bridge_in_reset.reset
			nios2_data_master_address                             => nios2_data_master_address,                                  --                               nios2_data_master.address
			nios2_data_master_waitrequest                         => nios2_data_master_waitrequest,                              --                                                .waitrequest
			nios2_data_master_byteenable                          => nios2_data_master_byteenable,                               --                                                .byteenable
			nios2_data_master_read                                => nios2_data_master_read,                                     --                                                .read
			nios2_data_master_readdata                            => nios2_data_master_readdata,                                 --                                                .readdata
			nios2_data_master_write                               => nios2_data_master_write,                                    --                                                .write
			nios2_data_master_writedata                           => nios2_data_master_writedata,                                --                                                .writedata
			nios2_data_master_debugaccess                         => nios2_data_master_debugaccess,                              --                                                .debugaccess
			nios2_instruction_master_address                      => nios2_instruction_master_address,                           --                        nios2_instruction_master.address
			nios2_instruction_master_waitrequest                  => nios2_instruction_master_waitrequest,                       --                                                .waitrequest
			nios2_instruction_master_read                         => nios2_instruction_master_read,                              --                                                .read
			nios2_instruction_master_readdata                     => nios2_instruction_master_readdata,                          --                                                .readdata
			nios2_debug_mem_slave_address                         => mm_interconnect_0_nios2_debug_mem_slave_address,            --                           nios2_debug_mem_slave.address
			nios2_debug_mem_slave_write                           => mm_interconnect_0_nios2_debug_mem_slave_write,              --                                                .write
			nios2_debug_mem_slave_read                            => mm_interconnect_0_nios2_debug_mem_slave_read,               --                                                .read
			nios2_debug_mem_slave_readdata                        => mm_interconnect_0_nios2_debug_mem_slave_readdata,           --                                                .readdata
			nios2_debug_mem_slave_writedata                       => mm_interconnect_0_nios2_debug_mem_slave_writedata,          --                                                .writedata
			nios2_debug_mem_slave_byteenable                      => mm_interconnect_0_nios2_debug_mem_slave_byteenable,         --                                                .byteenable
			nios2_debug_mem_slave_waitrequest                     => mm_interconnect_0_nios2_debug_mem_slave_waitrequest,        --                                                .waitrequest
			nios2_debug_mem_slave_debugaccess                     => mm_interconnect_0_nios2_debug_mem_slave_debugaccess,        --                                                .debugaccess
			onchip_flash_csr_address                              => mm_interconnect_0_onchip_flash_csr_address,                 --                                onchip_flash_csr.address
			onchip_flash_csr_write                                => mm_interconnect_0_onchip_flash_csr_write,                   --                                                .write
			onchip_flash_csr_read                                 => mm_interconnect_0_onchip_flash_csr_read,                    --                                                .read
			onchip_flash_csr_readdata                             => mm_interconnect_0_onchip_flash_csr_readdata,                --                                                .readdata
			onchip_flash_csr_writedata                            => mm_interconnect_0_onchip_flash_csr_writedata,               --                                                .writedata
			onchip_flash_data_address                             => mm_interconnect_0_onchip_flash_data_address,                --                               onchip_flash_data.address
			onchip_flash_data_write                               => mm_interconnect_0_onchip_flash_data_write,                  --                                                .write
			onchip_flash_data_read                                => mm_interconnect_0_onchip_flash_data_read,                   --                                                .read
			onchip_flash_data_readdata                            => mm_interconnect_0_onchip_flash_data_readdata,               --                                                .readdata
			onchip_flash_data_writedata                           => mm_interconnect_0_onchip_flash_data_writedata,              --                                                .writedata
			onchip_flash_data_burstcount                          => mm_interconnect_0_onchip_flash_data_burstcount,             --                                                .burstcount
			onchip_flash_data_readdatavalid                       => mm_interconnect_0_onchip_flash_data_readdatavalid,          --                                                .readdatavalid
			onchip_flash_data_waitrequest                         => mm_interconnect_0_onchip_flash_data_waitrequest,            --                                                .waitrequest
			onchip_ram_s1_address                                 => mm_interconnect_0_onchip_ram_s1_address,                    --                                   onchip_ram_s1.address
			onchip_ram_s1_write                                   => mm_interconnect_0_onchip_ram_s1_write,                      --                                                .write
			onchip_ram_s1_readdata                                => mm_interconnect_0_onchip_ram_s1_readdata,                   --                                                .readdata
			onchip_ram_s1_writedata                               => mm_interconnect_0_onchip_ram_s1_writedata,                  --                                                .writedata
			onchip_ram_s1_byteenable                              => mm_interconnect_0_onchip_ram_s1_byteenable,                 --                                                .byteenable
			onchip_ram_s1_chipselect                              => mm_interconnect_0_onchip_ram_s1_chipselect,                 --                                                .chipselect
			onchip_ram_s1_clken                                   => mm_interconnect_0_onchip_ram_s1_clken,                      --                                                .clken
			pio_led_s1_address                                    => mm_interconnect_0_pio_led_s1_address,                       --                                      pio_led_s1.address
			pio_led_s1_write                                      => mm_interconnect_0_pio_led_s1_write,                         --                                                .write
			pio_led_s1_readdata                                   => mm_interconnect_0_pio_led_s1_readdata,                      --                                                .readdata
			pio_led_s1_writedata                                  => mm_interconnect_0_pio_led_s1_writedata,                     --                                                .writedata
			pio_led_s1_chipselect                                 => mm_interconnect_0_pio_led_s1_chipselect,                    --                                                .chipselect
			pio_mode_s1_address                                   => mm_interconnect_0_pio_mode_s1_address,                      --                                     pio_mode_s1.address
			pio_mode_s1_readdata                                  => mm_interconnect_0_pio_mode_s1_readdata,                     --                                                .readdata
			pll_pll_slave_address                                 => mm_interconnect_0_pll_pll_slave_address,                    --                                   pll_pll_slave.address
			pll_pll_slave_write                                   => mm_interconnect_0_pll_pll_slave_write,                      --                                                .write
			pll_pll_slave_read                                    => mm_interconnect_0_pll_pll_slave_read,                       --                                                .read
			pll_pll_slave_readdata                                => mm_interconnect_0_pll_pll_slave_readdata,                   --                                                .readdata
			pll_pll_slave_writedata                               => mm_interconnect_0_pll_pll_slave_writedata,                  --                                                .writedata
			sdram_controller_s1_address                           => mm_interconnect_0_sdram_controller_s1_address,              --                             sdram_controller_s1.address
			sdram_controller_s1_write                             => mm_interconnect_0_sdram_controller_s1_write,                --                                                .write
			sdram_controller_s1_read                              => mm_interconnect_0_sdram_controller_s1_read,                 --                                                .read
			sdram_controller_s1_readdata                          => mm_interconnect_0_sdram_controller_s1_readdata,             --                                                .readdata
			sdram_controller_s1_writedata                         => mm_interconnect_0_sdram_controller_s1_writedata,            --                                                .writedata
			sdram_controller_s1_byteenable                        => mm_interconnect_0_sdram_controller_s1_byteenable,           --                                                .byteenable
			sdram_controller_s1_readdatavalid                     => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --                                                .readdatavalid
			sdram_controller_s1_waitrequest                       => mm_interconnect_0_sdram_controller_s1_waitrequest,          --                                                .waitrequest
			sdram_controller_s1_chipselect                        => mm_interconnect_0_sdram_controller_s1_chipselect,           --                                                .chipselect
			spi_flash_spi_control_port_address                    => mm_interconnect_0_spi_flash_spi_control_port_address,       --                      spi_flash_spi_control_port.address
			spi_flash_spi_control_port_write                      => mm_interconnect_0_spi_flash_spi_control_port_write,         --                                                .write
			spi_flash_spi_control_port_read                       => mm_interconnect_0_spi_flash_spi_control_port_read,          --                                                .read
			spi_flash_spi_control_port_readdata                   => mm_interconnect_0_spi_flash_spi_control_port_readdata,      --                                                .readdata
			spi_flash_spi_control_port_writedata                  => mm_interconnect_0_spi_flash_spi_control_port_writedata,     --                                                .writedata
			spi_flash_spi_control_port_chipselect                 => mm_interconnect_0_spi_flash_spi_control_port_chipselect,    --                                                .chipselect
			spi_g_sensor_spi_control_port_address                 => mm_interconnect_0_spi_g_sensor_spi_control_port_address,    --                   spi_g_sensor_spi_control_port.address
			spi_g_sensor_spi_control_port_write                   => mm_interconnect_0_spi_g_sensor_spi_control_port_write,      --                                                .write
			spi_g_sensor_spi_control_port_read                    => mm_interconnect_0_spi_g_sensor_spi_control_port_read,       --                                                .read
			spi_g_sensor_spi_control_port_readdata                => mm_interconnect_0_spi_g_sensor_spi_control_port_readdata,   --                                                .readdata
			spi_g_sensor_spi_control_port_writedata               => mm_interconnect_0_spi_g_sensor_spi_control_port_writedata,  --                                                .writedata
			spi_g_sensor_spi_control_port_chipselect              => mm_interconnect_0_spi_g_sensor_spi_control_port_chipselect, --                                                .chipselect
			sysid_control_slave_address                           => mm_interconnect_0_sysid_control_slave_address,              --                             sysid_control_slave.address
			sysid_control_slave_readdata                          => mm_interconnect_0_sysid_control_slave_readdata,             --                                                .readdata
			uart_s1_address                                       => mm_interconnect_0_uart_s1_address,                          --                                         uart_s1.address
			uart_s1_write                                         => mm_interconnect_0_uart_s1_write,                            --                                                .write
			uart_s1_read                                          => mm_interconnect_0_uart_s1_read,                             --                                                .read
			uart_s1_readdata                                      => mm_interconnect_0_uart_s1_readdata,                         --                                                .readdata
			uart_s1_writedata                                     => mm_interconnect_0_uart_s1_writedata,                        --                                                .writedata
			uart_s1_begintransfer                                 => mm_interconnect_0_uart_s1_begintransfer,                    --                                                .begintransfer
			uart_s1_chipselect                                    => mm_interconnect_0_uart_s1_chipselect                        --                                                .chipselect
		);

	irq_mapper : component NIOS_test_board_irq_mapper
		port map (
			clk           => pll_c0_clk,                     --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => nios2_irq_irq                   --    sender.irq
		);

	rst_controller : component nios_test_board_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios2_debug_reset_request_reset,    -- reset_in1.reset
			clk            => pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component nios_test_board_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios2_debug_reset_request_reset,    -- reset_in1.reset
			clk            => clk_in_clk,                         --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	mm_interconnect_0_pio_led_s1_write_ports_inv <= not mm_interconnect_0_pio_led_s1_write;

	mm_interconnect_0_uart_s1_read_ports_inv <= not mm_interconnect_0_uart_s1_read;

	mm_interconnect_0_uart_s1_write_ports_inv <= not mm_interconnect_0_uart_s1_write;

	mm_interconnect_0_spi_flash_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_flash_spi_control_port_read;

	mm_interconnect_0_spi_flash_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_flash_spi_control_port_write;

	mm_interconnect_0_spi_g_sensor_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_g_sensor_spi_control_port_read;

	mm_interconnect_0_spi_g_sensor_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_g_sensor_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of NIOS_test_board
